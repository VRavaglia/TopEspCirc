** Profile: "SCHEMATIC1-trans"  [ E:\ONEDRIVE - POLI.UFRJ.BR\MESTRADO\TOPESPCIRC\CompOrCad\Comp-PSpiceFiles\SCHEMATIC1\trans.sim ] 

** Creating circuit file "trans.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "C:\Cadence\SPB_16.5\tools\pspice\library\eval.lib" 
.lib "C:\Cadence\SPB_16.5\tools\pspice\library\CMOS35.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.3 0 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
